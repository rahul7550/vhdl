interface intf();
 logic sum;
 logic carry;
 logic a;
 logic b; 
endinterface
